/********** defines.v **********/
// `defines are only used to create type definitions (and in some local optimisations)
// module parameters should always be used locally in
// modules

`define OPT_MESHXYTURNS
`define DEBUG
`define X_ADDR_BITS 2
`define Y_ADDR_BITS 2
